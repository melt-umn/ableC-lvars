grammar edu:umn:cs:melt:exts:ableC:lvars:abstractsyntax;
