grammar edu:umn:cs:melt:exts:ableC:lvars;

exports edu:umn:cs:melt:exts:ableC:lvars:concretesyntax;
exports edu:umn:cs:melt:exts:ableC:lvars:abstractsyntax;
